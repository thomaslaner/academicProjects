library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.nes_controller_pkg.all;
use work.audio_cntrl_pkg.all;

package ball_game_pkg is

	type ball_game_state_t is (IDLE, PAUSED, RUNNING, GAME_OVER);


	component ball_game is
		generic (
			DISPLAY_WIDTH : integer;
			DISPLAY_HEIGHT : integer
		);
		port (
			clk : in std_logic;
			res_n : in std_logic;
			gfx_instr : out std_logic_vector(7 downto 0);
			gfx_instr_wr : out std_logic;
			gfx_instr_full : in std_logic;
			gfx_data : out std_logic_vector(15 downto 0);
			gfx_data_wr : out std_logic;
			gfx_data_full : in std_logic;
			gfx_frame_sync : in std_logic;
			controller : in nes_buttons_t;
			synth_cntrl : out synth_cntrl_vec_t(0 to 1);
			player_points : out std_logic_vector(15 downto 0);
			game_state : out ball_game_state_t
		);
	end component;

end package;

